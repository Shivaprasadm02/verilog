//--1--//
//diff bt monitor and strobe

//--2--//
//what is `timescale

//--3--//
//compiler directives and simulation directives

//--4--//
//how to write to a file

//--5--//
//explain $readmemb

//--6--//
//explain about $random

//--7--//
//limitations of timescale

//--8--//
"What is the display output for a, b?
module display_eg();
reg [2:0]a, b;
reg [2:0]c;
initial
begin
$strobe("1st a=%0d,b=%0d",a,b);
a='d4;
b='d7;
#10;
a='d6;
b='d2;
$strobe("2nd a=%0d,b=%0d",a,b);
#20;
b='d4;
a='d1;
end
endmodule"

//--9--//
"Explain the following Verilog code:
`timescale 10ns/100ps

module test;
reg [2:0]x;

initial
begin
#10.4567;
x=4;
end
endmodule"
//////

//--10--//
"Find the time-period of the below clk signal:
`timescale 1ns/1ns
reg clk;
initial
begin
#5 clk = 0;
forever #2.5 clk = ~clk;
end"
//time unit 2.5x1=2.5
//time period is 2.5x2=5 as precisoion is 1ns no fraction is allowed
//ans:-5ns

//-----------------11--------------////////////
What will be the output for the below snippet
`define MACRO1
`define MACRO2
module tb ( );
initial
begin
`ifdef MACRO1
$display (""This is MACRO1"");
`else
`ifdef MACRO2
$display (""This is MACRO2"");
`endif
`endif
end"
//ans:- This is MACRO1
//--12--//
What will be the time period of the clock (clk) generated by the following code segment?

`timescale 10ns/100ps
module test;
reg clk;
initial
#0.35 clk = 1’b0;
always #0.63 clk = ~clk;"
//0.63x10=6.3 and precision is 100ps=0.1ns so 6.3 is allowed
//timeperiod =6.3x2
//ans:- 12.6ns

//--13--//
Explain the below code?
reg clk;
integer count;
initial
begin
clk = 1'b0;
count = 0;
forever
#50 clk = ~clk;
end

always @ (posedge clk)
count = count + 1;

always @ (posedge clk)
$write (""count is equal to %d\n"", count)
//here its a race actually as we are reading before write
//evaluation of count are happening at 0time 
//if write was in same always block then it would have detected the change in value
//ans:- it displays previous value as write also starts at 0time 
//and assignmnet to count is not yet done when write executes

//--14--//
What is the hardware inferred from the below snippet?
always@(posedge clk or negedge reset)
begin
if(~reset)
b <= 1'b0;
else
begin
b <= a & b;
end
end
//synchronous ff with asynchronous clear
//ans:- it creates a dff with and gate as input

//--15--//
What is the hardware inferred from the below snippet?

always@(posedge clk1 or negedge clk2)
begin
if(~clk2 && a)
dout<=0;
else
dout<= din;
end
//a and din are sync to clk1
//not synthesizable
//ans:- 
//here clk2 is asynchronous and a is asynchronous,
//we cannot include both in an condition/expression

//--16--//
What are the values of A, B and C after the below code finishes executing?

reg [3:0] A, B, C;

initial
begin
$monitor(A,B,C);
A=0;
B=0;
C=0;
#1
A=B+1;
C=A+1;
B=C+1;
#1
A<=C+1;
C<=B+1;
B<=A+1;
end
//ans:-$monitor 
At 0ns : A=0 B=0 C =0
At 1ns : A=1 B=3 C =2
At 2ns : A=3 B=2 C =4

//--17--//
What logic is inferred by following snippet?

always@(posedge clk)
if(reset)
begin
c <= 0;
end
else if(s)
begin
c <=a;
end
//ans:- mux and ff

//--18--//
Whether the below snippet is valid code?

initial
begin
if( a )
MUX M1 (……);
else
DEC D1 (……) ;
end"

//--19--//
Predict the output of below snippet
always@(posedge clk or posedge rst)
if(rst)
x1= 0;
else
x1=x2;

always @ (posedge clk or posedge rst)
if ( rst )
x2 = 0;
else
x2 = x1;

//ans:- it creates a race condition

//--20--//
What is the value of r at 50ns?

reg [3:0] r;

initial
begin
r = 0;
r = #10 2;
r = #20 3;
#10;
r <= #20 4;
r <= #10 0;
end

//ans:- at 50 units 

///clock with 70% duty cycle
always
begin
clk = 1'b0;
#30;
clk = 1'b1;
#70;
end